interface up_if;
	logic up_clk;
	logic up_rst;
	logic[15:0] up_in;

	logic[15:0] up_out;
	logic up_eno;
	
endinterface: up_if