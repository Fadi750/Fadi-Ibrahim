interface relu_if;
	logic relu_clk;
	logic relu_reset;
	logic[19:0] relu_in;

	logic[19:0] relu_out;
	logic relu_en_o;
	
endinterface: relu_if