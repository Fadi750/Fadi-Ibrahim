module invsbox(datain,dataout);
  input [7:0] datain;
  output reg [7:0] dataout;
  
  always @(datain)
  begin
    case(datain)
  8'h00 :dataout= 8'h52;
  8'h01 :dataout= 8'h09;
  8'h02 :dataout= 8'h6a;
  8'h03 :dataout= 8'hd5;
  8'h04 :dataout= 8'h30;
  8'h05 :dataout= 8'h36;
  8'h06 :dataout= 8'ha5;
  8'h07 :dataout= 8'h38;
  8'h08 :dataout= 8'hbf;
  8'h09 :dataout= 8'h40;
  8'h0a :dataout= 8'ha3;
  8'h0b :dataout= 8'h9e;
  8'h0c :dataout= 8'h81;
  8'h0d :dataout= 8'hf3;
  8'h0e :dataout= 8'hd7;
  8'h0f :dataout= 8'hfb;
  8'h10 :dataout= 8'h7c;
  8'h11 :dataout= 8'he3;
  8'h12 :dataout= 8'h39;
  8'h13 :dataout= 8'h82;
  8'h14 :dataout= 8'h9b;
  8'h15 :dataout= 8'h2f;
  8'h16 :dataout= 8'hff;
  8'h17 :dataout= 8'h87;
  8'h18 :dataout= 8'h34;
  8'h19 :dataout= 8'h8e;
  8'h1a :dataout= 8'h43;
  8'h1b :dataout= 8'h44;
  8'h1c :dataout= 8'hc4;
  8'h1d :dataout= 8'hde;
  8'h1e :dataout= 8'he9;
  8'h1f :dataout= 8'hcb;
  8'h20 :dataout= 8'h54;
  8'h21 :dataout= 8'h7b;
  8'h22 :dataout= 8'h94;
  8'h23 :dataout= 8'h32;
  8'h24 :dataout= 8'ha6;
  8'h25 :dataout= 8'hc2;
  8'h26 :dataout= 8'h23;
  8'h27 :dataout= 8'h3d;
  8'h28 :dataout= 8'hee;
  8'h29 :dataout= 8'h4c;
  8'h2a :dataout= 8'h95;
  8'h2b :dataout= 8'h0b;
  8'h2c :dataout= 8'h42;
  8'h2d :dataout= 8'hfa;
  8'h2e :dataout= 8'hc3;
  8'h2f :dataout= 8'h4e;
  8'h30 :dataout= 8'h08;
  8'h31 :dataout= 8'h2e;
  8'h32 :dataout= 8'ha1;
  8'h33 :dataout= 8'h66;
  8'h34 :dataout= 8'h28;
  8'h35 :dataout= 8'hd9;
  8'h36 :dataout= 8'h24;
  8'h37 :dataout= 8'hb2;
  8'h38 :dataout= 8'h76;
  8'h39 :dataout= 8'h5b;
  8'h3a :dataout= 8'ha2;
  8'h3b :dataout= 8'h49;
  8'h3c :dataout= 8'h6d;
  8'h3d :dataout= 8'h8b;
  8'h3e :dataout= 8'hd1;
  8'h3f :dataout= 8'h25;
  8'h40 :dataout= 8'h72;
  8'h41 :dataout= 8'hf8;
  8'h42 :dataout= 8'hf6;
  8'h43 :dataout= 8'h64;
  8'h44 :dataout= 8'h86;
  8'h45 :dataout= 8'h68;
  8'h46 :dataout= 8'h98;
  8'h47 :dataout= 8'h16;
  8'h48 :dataout= 8'hd4;
  8'h49 :dataout= 8'ha4;
  8'h4a :dataout= 8'h5c;
  8'h4b :dataout= 8'hcc;
  8'h4c :dataout= 8'h5d;
  8'h4d :dataout= 8'h65;
  8'h4e :dataout= 8'hb6;
  8'h4f :dataout= 8'h92;
  8'h50 :dataout= 8'h6c;
  8'h51 :dataout= 8'h70;
  8'h52 :dataout= 8'h48;
  8'h53 :dataout= 8'h50;
  8'h54 :dataout= 8'hfd;
  8'h55 :dataout= 8'hed;
  8'h56 :dataout= 8'hb9;
  8'h57 :dataout= 8'hda;
  8'h58 :dataout= 8'h5e;
  8'h59 :dataout= 8'h15;
  8'h5a :dataout= 8'h46;
  8'h5b :dataout= 8'h57;
  8'h5c :dataout= 8'ha7;
  8'h5d :dataout= 8'h8d;
  8'h5e :dataout= 8'h9d;
  8'h5f :dataout= 8'h84;
  8'h60 :dataout= 8'h90;
  8'h61 :dataout= 8'hd8;
  8'h62 :dataout= 8'hab;
  8'h63 :dataout= 8'h00;
  8'h64 :dataout= 8'h8c;
  8'h65 :dataout= 8'hbc;
  8'h66 :dataout= 8'hd3;
  8'h67 :dataout= 8'h0a;
  8'h68 :dataout= 8'hf7;
  8'h69 :dataout= 8'he4;
  8'h6a :dataout= 8'h58;
  8'h6b :dataout= 8'h05;
  8'h6c :dataout= 8'hb8;
  8'h6d :dataout= 8'hb3;
  8'h6e :dataout= 8'h45;
  8'h6f :dataout= 8'h06;
  8'h70 :dataout= 8'hd0;
  8'h71 :dataout= 8'h2c;
  8'h72 :dataout= 8'h1e;
  8'h73 :dataout= 8'h8f;
  8'h74 :dataout= 8'hca;
  8'h75 :dataout= 8'h3f;
  8'h76 :dataout= 8'h0f;
  8'h77 :dataout= 8'h02;
  8'h78 :dataout= 8'hc1;
  8'h79 :dataout= 8'haf;
  8'h7a :dataout= 8'hbd;
  8'h7b :dataout= 8'h03;
  8'h7c :dataout= 8'h01;
  8'h7d :dataout= 8'h13;
  8'h7e :dataout= 8'h8a;
  8'h7f :dataout= 8'h6b;
  8'h80 :dataout= 8'h3a;
  8'h81 :dataout= 8'h91;
  8'h82 :dataout= 8'h11;
  8'h83 :dataout= 8'h41;
  8'h84 :dataout= 8'h4f;
  8'h85 :dataout= 8'h67;
  8'h86 :dataout= 8'hdc;
  8'h87 :dataout= 8'hea;
  8'h88 :dataout= 8'h97;
  8'h89 :dataout= 8'hf2;
  8'h8a :dataout= 8'hcf;
  8'h8b :dataout= 8'hce;
  8'h8c :dataout= 8'hf0;
  8'h8d :dataout= 8'hb4;
  8'h8e :dataout= 8'he6;
  8'h8f :dataout= 8'h73;
  8'h90 :dataout= 8'h96;
  8'h91 :dataout= 8'hac;
  8'h92 :dataout= 8'h74;
  8'h93 :dataout= 8'h22;
  8'h94 :dataout= 8'he7;
  8'h95 :dataout= 8'had;
  8'h96 :dataout= 8'h35;
  8'h97 :dataout= 8'h85;
  8'h98 :dataout= 8'he2;
  8'h99 :dataout= 8'hf9;
  8'h9a :dataout= 8'h37;
  8'h9b :dataout= 8'he8;
  8'h9c :dataout= 8'h1c;
  8'h9d :dataout= 8'h75;
  8'h9e :dataout= 8'hdf;
  8'h9f :dataout= 8'h6e;
  8'ha0 :dataout= 8'h47;
  8'ha1 :dataout= 8'hf1;
  8'ha2 :dataout= 8'h1a;
  8'ha3 :dataout= 8'h71;
  8'ha4 :dataout= 8'h1d;
  8'ha5 :dataout= 8'h29;
  8'ha6 :dataout= 8'hc5;
  8'ha7 :dataout= 8'h89;
  8'ha8 :dataout= 8'h6f;
  8'ha9 :dataout= 8'hb7;
  8'haa :dataout= 8'h62;
  8'hab :dataout= 8'h0e;
  8'hac :dataout= 8'haa;
  8'had :dataout= 8'h18;
  8'hae :dataout= 8'hbe;
  8'haf :dataout= 8'h1b;
  8'hb0 :dataout= 8'hfc;
  8'hb1 :dataout= 8'h56;
  8'hb2 :dataout= 8'h3e;
  8'hb3 :dataout= 8'h4b;
  8'hb4 :dataout= 8'hc6;
  8'hb5 :dataout= 8'hd2;
  8'hb6 :dataout= 8'h79;
  8'hb7 :dataout= 8'h20;
  8'hb8 :dataout= 8'h9a;
  8'hb9 :dataout= 8'hdb;
  8'hba :dataout= 8'hc0;
  8'hbb :dataout= 8'hfe;
  8'hbc :dataout= 8'h78;
  8'hbd :dataout= 8'hcd;
  8'hbe :dataout= 8'h5a;
  8'hbf :dataout= 8'hf4;
  8'hc0 :dataout= 8'h1f;
  8'hc1 :dataout= 8'hdd;
  8'hc2 :dataout= 8'ha8;
  8'hc3 :dataout= 8'h33;
  8'hc4 :dataout= 8'h88;
  8'hc5 :dataout= 8'h07;
  8'hc6 :dataout= 8'hc7;
  8'hc7 :dataout= 8'h31;
  8'hc8 :dataout= 8'hb1;
  8'hc9 :dataout= 8'h12;
  8'hca :dataout= 8'h10;
  8'hcb :dataout= 8'h59;
  8'hcc :dataout= 8'h27;
  8'hcd :dataout= 8'h80;
  8'hce :dataout= 8'hec;
  8'hcf :dataout= 8'h5f;
  8'hd0 :dataout= 8'h60;
  8'hd1 :dataout= 8'h51;
  8'hd2 :dataout= 8'h7f;
  8'hd3 :dataout= 8'ha9;
  8'hd4 :dataout= 8'h19;
  8'hd5 :dataout= 8'hb5;
  8'hd6 :dataout= 8'h4a;
  8'hd7 :dataout= 8'h0d;
  8'hd8 :dataout= 8'h2d;
  8'hd9 :dataout= 8'he5;
  8'hda :dataout= 8'h7a;
  8'hdb :dataout= 8'h9f;
  8'hdc :dataout= 8'h93;
  8'hdd :dataout= 8'hc9;
  8'hde :dataout= 8'h9c;
  8'hdf :dataout= 8'hef;
  8'he0 :dataout= 8'ha0;
  8'he1 :dataout= 8'he0;
  8'he2 :dataout= 8'h3b;
  8'he3 :dataout= 8'h4d;
  8'he4 :dataout= 8'hae;
  8'he5 :dataout= 8'h2a;
  8'he6 :dataout= 8'hf5;
  8'he7 :dataout= 8'hb0;
  8'he8 :dataout= 8'hc8;
  8'he9 :dataout= 8'heb;
  8'hea :dataout= 8'hbb;
  8'heb :dataout= 8'h3c;
  8'hec :dataout= 8'h83;
  8'hed :dataout= 8'h53;
  8'hee :dataout= 8'h99;
  8'hef :dataout= 8'h61;
  8'hf0 :dataout= 8'h17;
  8'hf1 :dataout= 8'h2b;
  8'hf2 :dataout= 8'h04;
  8'hf3 :dataout= 8'h7e;
  8'hf4 :dataout= 8'hba;
  8'hf5 :dataout= 8'h77;
  8'hf6 :dataout= 8'hd6;
  8'hf7 :dataout= 8'h26;
  8'hf8 :dataout= 8'he1;
  8'hf9 :dataout= 8'h69;
  8'hfa :dataout= 8'h14;
  8'hfb :dataout= 8'h63;
  8'hfc :dataout= 8'h55;
  8'hfd :dataout= 8'h21;
  8'hfe :dataout= 8'h0c;
  8'hff :dataout= 8'h7d;
endcase
end
endmodule

  