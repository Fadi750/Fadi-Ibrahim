package up_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "up_sequencer.svh"
	`include "up_driver.svh"
	`include "up_monitor.svh"
	`include "up_agent.svh"
	`include "up_scoreboard.svh"
	`include "up_env.svh"
	`include "up_test.svh"
	`include "up_config.svh"
	
endpackage: up_pkg