package relu_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "relu_sequencer.svh"
	`include "relu_driver.svh"
	`include "relu_monitor.svh"
	`include "relu_agent.svh"
	`include "relu_scoreboard.svh"
	`include "relu_env.svh"
	`include "relu_test.svh"
	`include "relu_config.svh"
	
endpackage: relu_pkg
