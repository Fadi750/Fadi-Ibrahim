package cvpu_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "cvpu_sequencer.svh"
	`include "cvpu_driver.svh"
	`include "cvpu_monitor.svh"
	`include "cvpu_agent.svh"
	`include "cvpu_scoreboard.svh"
	`include "cvpu_env.svh"
	`include "cvpu_test.svh"
	`include "cvpu_config.svh"
	
endpackage: cvpu_pkg