module inv_shift(s,ss);
  input [127:0] s;
  output reg [127:0] ss;
   
    
    always@(s) begin 
      ss[7:0]<=s[103:96];
      ss[15:8]<=s[79:72];
      ss[23:16]<=s[55:48];
      ss[31:24]<=s[31:24];
      ss[39:32]<=s[7:0];
      ss[47:40]<=s[111:104];
      ss[55:48]<=s[87:80];
      ss[63:56]<=s[63:56];
      ss[71:64]<=s[39:32];
      ss[79:72]<=s[15:8];
      ss[87:80]<=s[119:112];
      ss[95:88]<=s[95:88];
      ss[103:96]<=s[71:64];
      ss[111:104]<=s[47:40];
      ss[119:112]<=s[23:16];
      ss[127:120]<=s[127:120];
    end
  endmodule
